magic
tech scmos
timestamp 1636276523
<< nwell >>
rect -12 2 37 18
<< polysilicon >>
rect -20 14 10 16
rect -20 -14 -18 14
rect -8 10 -6 12
rect 8 10 10 14
rect 29 10 31 12
rect -8 -2 -6 4
rect 8 2 10 4
rect 29 2 31 4
rect 8 0 31 2
rect -8 -4 10 -2
rect -8 -8 -6 -6
rect 8 -8 10 -4
rect 29 -8 31 0
rect -8 -14 -6 -11
rect -20 -16 -6 -14
rect 8 -15 10 -11
rect 29 -13 31 -11
rect 8 -17 17 -15
<< ndiffusion >>
rect -9 -11 -8 -8
rect -6 -11 -5 -8
rect 7 -11 8 -8
rect 10 -11 11 -8
rect 28 -11 29 -8
rect 31 -11 32 -8
<< pdiffusion >>
rect -11 9 -8 10
rect -9 5 -8 9
rect -11 4 -8 5
rect -6 9 -3 10
rect 5 9 8 10
rect -6 5 -5 9
rect 7 5 8 9
rect -6 4 -3 5
rect 5 4 8 5
rect 10 9 13 10
rect 26 9 29 10
rect 10 5 11 9
rect 28 5 29 9
rect 10 4 13 5
rect 26 4 29 5
rect 31 9 34 10
rect 31 5 32 9
rect 31 4 34 5
<< metal1 >>
rect -4 18 15 21
rect -4 9 -1 18
rect 12 9 15 18
rect 25 14 32 17
rect 25 9 28 14
rect -13 -7 -10 5
rect -4 -7 -1 5
rect 3 -7 6 5
rect 12 -7 15 5
rect 33 -1 36 5
rect 18 -4 36 -1
rect 18 -14 21 -4
rect 33 -7 36 -4
rect 24 -15 27 -11
rect 24 -18 33 -15
<< ntransistor >>
rect -8 -11 -6 -8
rect 8 -11 10 -8
rect 29 -11 31 -8
<< ptransistor >>
rect -8 4 -6 10
rect 8 4 10 10
rect 29 4 31 10
<< polycontact >>
rect 17 -18 21 -14
<< ndcontact >>
rect -13 -11 -9 -7
rect -5 -11 -1 -7
rect 3 -11 7 -7
rect 11 -11 15 -7
rect 24 -11 28 -7
rect 32 -11 36 -7
<< pdcontact >>
rect -13 5 -9 9
rect -5 5 -1 9
rect 3 5 7 9
rect 11 5 15 9
rect 24 5 28 9
rect 32 5 36 9
<< psubstratepcontact >>
rect 33 -19 37 -15
<< nsubstratencontact >>
rect 32 14 36 18
<< labels >>
rlabel metal1 5 19 5 19 1 Out
rlabel metal1 29 -17 29 -17 1 Vss
rlabel metal1 30 15 30 15 1 Vdd
rlabel metal1 34 -3 34 -3 1 S_bar
rlabel polysilicon 30 1 30 1 1 S
rlabel metal1 4 0 4 0 3 I1
rlabel metal1 -12 0 -12 0 3 I0
rlabel polysilicon -19 0 -19 0 1 S
rlabel polysilicon -7 -3 -7 -3 1 S_bar
<< end >>
