* SPICE3 file created from nor2.ext - technology: scmos

.option scale=1u

M1000 out a vss Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 d1s2 a vdd w_n14_7# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out b d1s2 w_n14_7# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vss b out Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vss Gnd 4.51fF
C1 out Gnd 3.38fF
C2 b Gnd 5.71fF
C3 a Gnd 5.71fF
C4 vdd Gnd 2.68fF
