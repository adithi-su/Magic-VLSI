magic
tech scmos
timestamp 1636303986
<< nwell >>
rect 11 25 60 42
<< polysilicon >>
rect 16 33 18 35
rect 36 33 38 35
rect 52 33 54 35
rect 16 25 18 27
rect 17 21 18 25
rect 16 10 18 21
rect 36 18 38 27
rect 52 25 54 27
rect 53 21 54 25
rect 37 14 38 18
rect 36 10 38 14
rect 52 10 54 21
rect 16 5 18 7
rect 36 5 38 7
rect 52 4 54 7
<< ndiffusion >>
rect 15 7 16 10
rect 18 7 36 10
rect 38 7 39 10
rect 51 7 52 10
rect 54 7 55 10
<< pdiffusion >>
rect 13 32 16 33
rect 15 28 16 32
rect 13 27 16 28
rect 18 32 21 33
rect 33 32 36 33
rect 18 28 19 32
rect 35 28 36 32
rect 18 27 21 28
rect 33 27 36 28
rect 38 32 41 33
rect 48 32 52 33
rect 38 28 39 32
rect 51 28 52 32
rect 38 27 41 28
rect 48 27 52 28
rect 54 32 58 33
rect 54 28 56 32
rect 54 27 58 28
<< metal1 >>
rect 15 38 31 41
rect 35 38 47 41
rect 12 32 15 38
rect 31 32 34 38
rect 47 32 50 38
rect 20 25 23 28
rect 40 25 43 28
rect 20 22 49 25
rect 40 11 43 22
rect 56 11 59 28
rect 11 3 14 7
rect 47 3 50 7
rect 15 -1 46 2
<< ntransistor >>
rect 16 7 18 10
rect 36 7 38 10
rect 52 7 54 10
<< ptransistor >>
rect 16 27 18 33
rect 36 27 38 33
rect 52 27 54 33
<< polycontact >>
rect 13 21 17 25
rect 49 21 53 25
rect 33 14 37 18
<< ndcontact >>
rect 11 7 15 11
rect 39 7 43 11
rect 47 7 51 11
rect 55 7 59 11
<< pdcontact >>
rect 11 28 15 32
rect 19 28 23 32
rect 31 28 35 32
rect 39 28 43 32
rect 47 28 51 32
rect 56 28 60 32
<< psubstratepcontact >>
rect 11 -1 15 3
rect 46 -1 50 3
<< nsubstratencontact >>
rect 11 38 15 42
rect 31 38 35 42
rect 47 38 51 42
<< labels >>
rlabel metal1 22 39 22 39 1 Vdd
rlabel metal1 22 0 22 0 1 Gnd
rlabel metal1 57 18 57 18 3 Out
<< end >>
