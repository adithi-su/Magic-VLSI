* SPICE3 file created from nor3.ext - technology: scmos

.option scale=1u

M1000 d1s2 A vdd vdd pfet w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 d2s3 B d1s2 vdd pfet w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out C vss Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vss B out Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 out C d2s3 vdd pfet w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out A vss Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vss Gnd 3.85fF
C1 out Gnd 4.79fF
C2 C Gnd 5.47fF
C3 B Gnd 5.47fF
C4 A Gnd 5.47fF
