* SPICE3 file created from HA.ext - technology: scmos

.option scale=1u

M1000 a_75_28# in Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 in B Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_75_77# in a_75_57# Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_75_77# A Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 sum a_75_28# a_133_47# Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 sum a_75_77# Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_13_34# A Gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_75_28# B Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 carry in Gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_75_77# in Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 sum a_75_28# Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 in B a_13_34# Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 in A Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 a_75_57# A Gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 a_75_28# B a_75_8# Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 a_133_47# a_75_77# Gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 a_75_8# in Gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 carry in Vdd Vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 Vdd A 4.15fF
C1 Vdd B 2.86fF
C2 Vdd a_75_77# 2.42fF
C3 Vdd in 5.46fF
C4 Vdd a_75_28# 2.18fF
C5 sum Gnd 4.51fF
C6 a_75_28# Gnd 20.84fF
C7 Gnd Gnd 33.16fF
C8 B Gnd 30.27fF
C9 a_75_77# Gnd 13.69fF
C10 in Gnd 44.15fF
C11 A Gnd 24.29fF
C12 Vdd Gnd 30.04fF
