magic
tech scmos
timestamp 1636295556
<< nwell >>
rect -79 154 -62 186
rect 21 134 37 183
rect -105 92 -88 124
rect -56 92 -39 124
rect -78 34 -61 66
rect -79 -13 -62 19
rect -105 -75 -88 -43
rect -56 -75 -39 -43
rect -78 -133 -61 -101
<< polysilicon >>
rect 3 189 12 191
rect 16 189 35 191
rect -99 179 -97 181
rect -94 180 -83 181
rect -79 180 -77 181
rect -94 179 -77 180
rect -71 179 -69 181
rect 3 179 5 189
rect 3 177 8 179
rect 11 177 13 179
rect 15 177 23 179
rect 29 177 31 179
rect -99 159 -97 161
rect -94 160 -90 161
rect 15 163 17 177
rect 33 163 35 189
rect 2 161 8 163
rect 11 161 17 163
rect 19 161 23 163
rect 29 161 35 163
rect -86 160 -77 161
rect -94 159 -77 160
rect -71 159 -69 161
rect 2 154 4 161
rect 19 142 21 161
rect 6 140 8 142
rect 11 140 23 142
rect 29 140 31 142
rect -125 117 -123 119
rect -120 118 -109 119
rect -105 118 -103 119
rect -120 117 -103 118
rect -97 117 -95 119
rect -76 117 -74 119
rect -71 118 -60 119
rect -56 118 -54 119
rect -71 117 -54 118
rect -48 117 -46 119
rect -125 97 -123 99
rect -120 98 -116 99
rect -112 98 -103 99
rect -120 97 -103 98
rect -97 97 -95 99
rect -76 97 -74 99
rect -71 98 -67 99
rect -63 98 -54 99
rect -71 97 -54 98
rect -48 97 -46 99
rect -98 59 -96 61
rect -93 60 -82 61
rect -78 60 -76 61
rect -93 59 -76 60
rect -70 59 -68 61
rect -98 39 -96 41
rect -93 40 -89 41
rect -85 40 -76 41
rect -93 39 -76 40
rect -70 39 -68 41
rect -99 12 -97 14
rect -94 13 -83 14
rect -79 13 -77 14
rect -94 12 -77 13
rect -71 12 -69 14
rect -99 -8 -97 -6
rect -94 -7 -90 -6
rect -86 -7 -77 -6
rect -94 -8 -77 -7
rect -71 -8 -69 -6
rect -125 -50 -123 -48
rect -120 -49 -109 -48
rect -105 -49 -103 -48
rect -120 -50 -103 -49
rect -97 -50 -95 -48
rect -76 -50 -74 -48
rect -71 -49 -60 -48
rect -56 -49 -54 -48
rect -71 -50 -54 -49
rect -48 -50 -46 -48
rect -125 -70 -123 -68
rect -120 -69 -116 -68
rect -112 -69 -103 -68
rect -120 -70 -103 -69
rect -97 -70 -95 -68
rect -76 -70 -74 -68
rect -71 -69 -67 -68
rect -63 -69 -54 -68
rect -71 -70 -54 -69
rect -48 -70 -46 -68
rect -98 -108 -96 -106
rect -93 -107 -82 -106
rect -78 -107 -76 -106
rect -93 -108 -76 -107
rect -70 -108 -68 -106
rect -98 -128 -96 -126
rect -93 -127 -89 -126
rect -85 -127 -76 -126
rect -93 -128 -76 -127
rect -70 -128 -68 -126
<< ndiffusion >>
rect -97 181 -94 182
rect 8 179 11 180
rect -97 161 -94 179
rect 8 176 11 177
rect 8 163 11 164
rect -97 158 -94 159
rect 8 160 11 161
rect 8 142 11 143
rect 8 139 11 140
rect -123 119 -120 120
rect -74 119 -71 120
rect -123 99 -120 117
rect -74 99 -71 117
rect -123 96 -120 97
rect -74 96 -71 97
rect -96 61 -93 62
rect -96 41 -93 59
rect -96 38 -93 39
rect -97 14 -94 15
rect -97 -6 -94 12
rect -97 -9 -94 -8
rect -123 -48 -120 -47
rect -74 -48 -71 -47
rect -123 -68 -120 -50
rect -74 -68 -71 -50
rect -123 -71 -120 -70
rect -74 -71 -71 -70
rect -96 -106 -93 -105
rect -96 -126 -93 -108
rect -96 -129 -93 -128
<< pdiffusion >>
rect -77 182 -76 184
rect -72 182 -71 184
rect -77 181 -71 182
rect 23 180 24 182
rect 28 180 29 182
rect 23 179 29 180
rect -77 178 -71 179
rect -77 176 -76 178
rect -72 176 -71 178
rect -77 162 -76 164
rect -72 162 -71 164
rect 23 176 29 177
rect 23 174 24 176
rect 28 174 29 176
rect 23 164 24 166
rect 28 164 29 166
rect 23 163 29 164
rect -77 161 -71 162
rect -77 158 -71 159
rect -77 156 -76 158
rect -72 156 -71 158
rect 23 160 29 161
rect 23 158 24 160
rect 28 158 29 160
rect 23 143 24 145
rect 28 143 29 145
rect 23 142 29 143
rect 23 139 29 140
rect 23 137 24 139
rect 28 137 29 139
rect -103 120 -102 122
rect -98 120 -97 122
rect -103 119 -97 120
rect -54 120 -53 122
rect -49 120 -48 122
rect -54 119 -48 120
rect -103 116 -97 117
rect -103 114 -102 116
rect -98 114 -97 116
rect -103 100 -102 102
rect -98 100 -97 102
rect -103 99 -97 100
rect -54 116 -48 117
rect -54 114 -53 116
rect -49 114 -48 116
rect -54 100 -53 102
rect -49 100 -48 102
rect -54 99 -48 100
rect -103 96 -97 97
rect -103 94 -102 96
rect -98 94 -97 96
rect -54 96 -48 97
rect -54 94 -53 96
rect -49 94 -48 96
rect -76 62 -75 64
rect -71 62 -70 64
rect -76 61 -70 62
rect -76 58 -70 59
rect -76 56 -75 58
rect -71 56 -70 58
rect -76 42 -75 44
rect -71 42 -70 44
rect -76 41 -70 42
rect -76 38 -70 39
rect -76 36 -75 38
rect -71 36 -70 38
rect -77 15 -76 17
rect -72 15 -71 17
rect -77 14 -71 15
rect -77 11 -71 12
rect -77 9 -76 11
rect -72 9 -71 11
rect -77 -5 -76 -3
rect -72 -5 -71 -3
rect -77 -6 -71 -5
rect -77 -9 -71 -8
rect -77 -11 -76 -9
rect -72 -11 -71 -9
rect -103 -47 -102 -45
rect -98 -47 -97 -45
rect -103 -48 -97 -47
rect -54 -47 -53 -45
rect -49 -47 -48 -45
rect -54 -48 -48 -47
rect -103 -51 -97 -50
rect -103 -53 -102 -51
rect -98 -53 -97 -51
rect -103 -67 -102 -65
rect -98 -67 -97 -65
rect -103 -68 -97 -67
rect -54 -51 -48 -50
rect -54 -53 -53 -51
rect -49 -53 -48 -51
rect -54 -67 -53 -65
rect -49 -67 -48 -65
rect -54 -68 -48 -67
rect -103 -71 -97 -70
rect -103 -73 -102 -71
rect -98 -73 -97 -71
rect -54 -71 -48 -70
rect -54 -73 -53 -71
rect -49 -73 -48 -71
rect -76 -105 -75 -103
rect -71 -105 -70 -103
rect -76 -106 -70 -105
rect -76 -109 -70 -108
rect -76 -111 -75 -109
rect -71 -111 -70 -109
rect -76 -125 -75 -123
rect -71 -125 -70 -123
rect -76 -126 -70 -125
rect -76 -129 -70 -128
rect -76 -131 -75 -129
rect -71 -131 -70 -129
<< metal1 >>
rect -115 190 -103 192
rect 13 193 16 198
rect -99 190 -86 192
rect -115 189 -86 190
rect -130 164 -127 182
rect -130 138 -127 160
rect -130 124 -127 134
rect -127 121 -123 124
rect -130 96 -127 120
rect -115 102 -112 189
rect -105 183 -97 186
rect -89 164 -86 189
rect -82 189 -71 192
rect -67 189 -56 192
rect -82 184 -79 189
rect -72 182 -66 185
rect -59 184 -56 189
rect -82 174 -76 177
rect -66 176 -63 182
rect -59 181 8 184
rect -82 157 -79 174
rect -66 166 -63 172
rect -72 163 -66 166
rect -93 154 -76 157
rect -82 148 -79 154
rect -108 145 -64 148
rect -108 122 -105 145
rect -92 124 -89 128
rect -82 124 -79 135
rect -98 120 -92 123
rect -78 121 -74 124
rect -108 112 -102 115
rect -108 95 -105 112
rect -92 104 -89 120
rect -98 101 -92 104
rect -67 102 -64 145
rect -59 122 -56 181
rect 12 181 24 184
rect 12 172 24 175
rect 28 172 40 175
rect -43 132 -40 172
rect 37 169 40 172
rect -22 165 8 168
rect -43 124 -40 128
rect -49 120 -43 123
rect -43 116 -40 120
rect -59 112 -53 115
rect -119 92 -102 95
rect -59 95 -56 112
rect -43 104 -40 112
rect -49 101 -43 104
rect -70 92 -53 95
rect -130 67 -127 92
rect -108 89 -105 92
rect -67 89 -64 92
rect -108 86 -86 89
rect -127 63 -104 66
rect -130 19 -127 63
rect -100 63 -96 66
rect -89 44 -86 86
rect -81 86 -64 89
rect -81 64 -78 86
rect -43 66 -40 100
rect -71 62 -65 65
rect -61 62 -43 65
rect -81 54 -75 57
rect -81 37 -78 54
rect -65 46 -62 62
rect -71 43 -65 46
rect -92 34 -75 37
rect -89 31 -86 34
rect -22 31 -19 165
rect 12 165 24 168
rect 37 165 39 169
rect 12 156 24 159
rect 37 159 40 165
rect 28 156 40 159
rect 5 150 18 153
rect 1 144 8 147
rect 1 138 4 144
rect -10 135 0 138
rect 15 138 18 150
rect 28 143 36 146
rect 33 139 36 143
rect 12 135 24 138
rect 33 115 36 135
rect -89 28 -19 31
rect -89 25 -86 28
rect -130 -3 -127 15
rect -130 -29 -127 -7
rect -130 -43 -127 -33
rect -115 22 -86 25
rect -127 -46 -123 -43
rect -130 -71 -127 -47
rect -115 -65 -112 22
rect -105 16 -97 19
rect -89 -3 -86 22
rect -82 22 -56 25
rect -82 17 -79 22
rect -72 15 -66 18
rect -82 7 -76 10
rect -66 9 -63 15
rect -82 -10 -79 7
rect -66 -1 -63 5
rect -72 -4 -66 -1
rect -93 -13 -76 -10
rect -82 -19 -79 -13
rect -108 -22 -64 -19
rect -108 -45 -105 -22
rect -92 -43 -89 -39
rect -82 -43 -79 -32
rect -98 -47 -92 -44
rect -78 -46 -74 -43
rect -108 -55 -102 -52
rect -108 -72 -105 -55
rect -92 -63 -89 -47
rect -98 -66 -92 -63
rect -67 -65 -64 -22
rect -59 -45 -56 22
rect -43 -35 -40 5
rect -43 -43 -40 -39
rect -49 -47 -43 -44
rect -59 -55 -53 -52
rect -119 -75 -102 -72
rect -59 -72 -56 -55
rect -43 -63 -40 -47
rect -49 -66 -43 -63
rect -70 -75 -53 -72
rect -130 -100 -127 -75
rect -108 -78 -105 -75
rect -67 -78 -64 -75
rect -108 -81 -86 -78
rect -127 -104 -104 -101
rect -100 -104 -96 -101
rect -89 -123 -86 -81
rect -81 -81 -64 -78
rect -81 -103 -78 -81
rect -43 -101 -40 -67
rect -71 -105 -65 -102
rect -61 -105 -43 -102
rect -81 -113 -75 -110
rect -81 -130 -78 -113
rect -65 -121 -62 -105
rect -71 -124 -65 -121
rect -92 -133 -85 -130
rect -81 -133 -75 -130
<< metal2 >>
rect -102 194 -99 198
rect -70 193 -67 198
rect -127 183 -109 186
rect -62 172 -43 175
rect 43 166 47 169
rect -130 138 -82 139
rect -127 136 -82 138
rect -78 136 -14 139
rect -88 128 -43 131
rect -39 112 32 115
rect -127 16 -109 19
rect -43 9 -40 63
rect -62 5 -43 8
rect -130 -29 -82 -28
rect -127 -31 -82 -29
rect -88 -39 -43 -36
rect -84 -139 -81 -134
<< ntransistor >>
rect -97 179 -94 181
rect 8 177 11 179
rect -97 159 -94 161
rect 8 161 11 163
rect 8 140 11 142
rect -123 117 -120 119
rect -74 117 -71 119
rect -123 97 -120 99
rect -74 97 -71 99
rect -96 59 -93 61
rect -96 39 -93 41
rect -97 12 -94 14
rect -97 -8 -94 -6
rect -123 -50 -120 -48
rect -74 -50 -71 -48
rect -123 -70 -120 -68
rect -74 -70 -71 -68
rect -96 -108 -93 -106
rect -96 -128 -93 -126
<< ptransistor >>
rect -77 179 -71 181
rect 23 177 29 179
rect 23 161 29 163
rect -77 159 -71 161
rect 23 140 29 142
rect -103 117 -97 119
rect -54 117 -48 119
rect -103 97 -97 99
rect -54 97 -48 99
rect -76 59 -70 61
rect -76 39 -70 41
rect -77 12 -71 14
rect -77 -8 -71 -6
rect -103 -50 -97 -48
rect -54 -50 -48 -48
rect -103 -70 -97 -68
rect -54 -70 -48 -68
rect -76 -108 -70 -106
rect -76 -128 -70 -126
<< polycontact >>
rect 12 189 16 193
rect -83 180 -79 184
rect -90 160 -86 164
rect 1 150 5 154
rect -109 118 -105 122
rect -60 118 -56 122
rect -116 98 -112 102
rect -67 98 -63 102
rect -82 60 -78 64
rect -89 40 -85 44
rect -83 13 -79 17
rect -90 -7 -86 -3
rect -109 -49 -105 -45
rect -60 -49 -56 -45
rect -116 -69 -112 -65
rect -67 -69 -63 -65
rect -82 -107 -78 -103
rect -89 -127 -85 -123
<< ndcontact >>
rect -97 182 -93 186
rect 8 180 12 184
rect 8 172 12 176
rect 8 164 12 168
rect -97 154 -93 158
rect 8 156 12 160
rect 8 143 12 147
rect 8 135 12 139
rect -123 120 -119 124
rect -74 120 -70 124
rect -123 92 -119 96
rect -74 92 -70 96
rect -96 62 -92 66
rect -96 34 -92 38
rect -97 15 -93 19
rect -97 -13 -93 -9
rect -123 -47 -119 -43
rect -74 -47 -70 -43
rect -123 -75 -119 -71
rect -74 -75 -70 -71
rect -96 -105 -92 -101
rect -96 -133 -92 -129
<< pdcontact >>
rect -76 182 -72 186
rect 24 180 28 184
rect -76 174 -72 178
rect -76 162 -72 166
rect 24 172 28 176
rect 24 164 28 168
rect -76 154 -72 158
rect 24 156 28 160
rect 24 143 28 147
rect 24 135 28 139
rect -102 120 -98 124
rect -53 120 -49 124
rect -102 112 -98 116
rect -102 100 -98 104
rect -53 112 -49 116
rect -53 100 -49 104
rect -102 92 -98 96
rect -53 92 -49 96
rect -75 62 -71 66
rect -75 54 -71 58
rect -75 42 -71 46
rect -75 34 -71 38
rect -76 15 -72 19
rect -76 7 -72 11
rect -76 -5 -72 -1
rect -76 -13 -72 -9
rect -102 -47 -98 -43
rect -53 -47 -49 -43
rect -102 -55 -98 -51
rect -102 -67 -98 -63
rect -53 -55 -49 -51
rect -53 -67 -49 -63
rect -102 -75 -98 -71
rect -53 -75 -49 -71
rect -75 -105 -71 -101
rect -75 -113 -71 -109
rect -75 -125 -71 -121
rect -75 -133 -71 -129
<< m2contact >>
rect -103 190 -99 194
rect -131 182 -127 186
rect -131 134 -127 138
rect -109 182 -105 186
rect -71 189 -67 193
rect -66 172 -62 176
rect -82 135 -78 139
rect -92 128 -88 132
rect -43 172 -39 176
rect -43 128 -39 132
rect -43 112 -39 116
rect 39 165 43 169
rect -14 135 -10 139
rect 32 111 36 115
rect -131 15 -127 19
rect -131 -33 -127 -29
rect -109 15 -105 19
rect -66 5 -62 9
rect -82 -32 -78 -28
rect -92 -39 -88 -35
rect -43 5 -39 9
rect -43 -39 -39 -35
rect -85 -134 -81 -130
<< psubstratepcontact >>
rect -131 160 -127 164
rect 0 134 4 138
rect -131 120 -127 124
rect -82 120 -78 124
rect -131 92 -127 96
rect -131 63 -127 67
rect -104 62 -100 66
rect -131 -7 -127 -3
rect -131 -47 -127 -43
rect -82 -47 -78 -43
rect -131 -75 -127 -71
rect -131 -104 -127 -100
rect -104 -105 -100 -101
<< nsubstratencontact >>
rect -66 182 -62 186
rect -66 162 -62 166
rect 33 135 37 139
rect -92 120 -88 124
rect -43 120 -39 124
rect -92 100 -88 104
rect -43 100 -39 104
rect -65 62 -61 66
rect -43 62 -39 66
rect -65 42 -61 46
rect -66 15 -62 19
rect -66 -5 -62 -1
rect -92 -47 -88 -43
rect -43 -47 -39 -43
rect -92 -67 -88 -63
rect -43 -67 -39 -63
rect -65 -105 -61 -101
rect -43 -105 -39 -101
rect -65 -125 -61 -121
<< labels >>
rlabel metal1 -114 24 -114 24 3 B
rlabel metal1 -129 -13 -129 -13 3 Gnd
rlabel metal1 -42 -16 -42 -16 3 Vdd
rlabel metal1 -58 191 -58 191 3 A
rlabel polycontact -58 120 -58 120 3 A
rlabel polycontact -81 182 -81 182 3 A
rlabel polycontact -114 100 -114 100 3 B
rlabel polycontact -88 162 -88 162 3 B
rlabel metal1 -114 191 -114 191 3 B
rlabel metal1 -129 154 -129 154 3 Gnd
rlabel metal1 -42 151 -42 151 3 Vdd
rlabel polycontact -81 15 -81 15 1 A2
rlabel polycontact -88 -5 -88 -5 1 B2
rlabel metal1 -58 24 -58 24 5 A2
rlabel polycontact -58 -47 -58 -47 1 A2
rlabel polycontact -114 -67 -114 -67 1 B2
rlabel metal1 -88 35 -88 35 1 Out1
rlabel m2contact -83 -132 -83 -132 1 sum
rlabel polysilicon 16 178 16 178 3 S_bar
rlabel polysilicon 19 190 19 190 3 S
rlabel metal1 19 183 19 183 5 I0
rlabel metal1 19 167 19 167 5 I1
rlabel polysilicon 20 141 20 141 3 S
rlabel metal1 16 137 16 137 3 S_bar
rlabel metal1 34 141 34 141 3 Vdd
rlabel metal2 45 167 45 167 1 carry
rlabel metal1 14 195 14 195 1 Ci
rlabel metal2 -69 196 -69 196 1 A
rlabel metal2 -101 196 -101 196 1 B
rlabel metal1 2 142 2 142 1 Gnd
<< end >>
