magic
tech scmos
timestamp 1635711947
<< nwell >>
rect 0 31 43 49
<< polysilicon >>
rect 7 40 9 42
rect 18 40 20 42
rect 35 40 37 42
rect 7 28 9 34
rect 18 30 20 34
rect 8 24 9 28
rect 19 26 20 30
rect 7 16 9 24
rect 18 16 20 26
rect 35 24 37 34
rect 36 20 37 24
rect 35 16 37 20
rect 7 7 9 10
rect 18 7 20 10
rect 35 7 37 10
<< ndiffusion >>
rect 2 15 7 16
rect 5 11 7 15
rect 2 10 7 11
rect 9 15 18 16
rect 9 11 12 15
rect 16 11 18 15
rect 9 10 18 11
rect 20 15 35 16
rect 20 11 22 15
rect 26 11 35 15
rect 20 10 35 11
rect 37 15 42 16
rect 37 11 40 15
rect 37 10 42 11
<< pdiffusion >>
rect 2 39 7 40
rect 5 35 7 39
rect 2 34 7 35
rect 9 34 18 40
rect 20 39 35 40
rect 20 35 22 39
rect 26 35 29 39
rect 33 35 35 39
rect 20 34 35 35
rect 37 39 42 40
rect 37 35 40 39
rect 37 34 42 35
<< metal1 >>
rect 1 46 14 49
rect 18 46 32 49
rect 1 39 4 46
rect 29 39 32 46
rect 23 23 26 35
rect 12 20 32 23
rect 12 15 15 20
rect 40 15 43 35
rect 2 5 5 11
rect 23 5 26 11
rect 2 4 26 5
rect 2 2 13 4
rect 17 2 26 4
<< ntransistor >>
rect 7 10 9 16
rect 18 10 20 16
rect 35 10 37 16
<< ptransistor >>
rect 7 34 9 40
rect 18 34 20 40
rect 35 34 37 40
<< polycontact >>
rect 4 24 8 28
rect 15 26 19 30
rect 32 20 36 24
<< ndcontact >>
rect 1 11 5 15
rect 12 11 16 15
rect 22 11 26 15
rect 40 11 44 15
<< pdcontact >>
rect 1 35 5 39
rect 22 35 26 39
rect 29 35 33 39
rect 40 35 44 39
<< psubstratepcontact >>
rect 13 0 17 4
<< nsubstratencontact >>
rect 14 46 18 50
<< labels >>
rlabel metal1 9 47 9 47 1 vdd
rlabel metal1 8 3 8 3 1 vss
rlabel polycontact 6 26 6 26 1 a
rlabel polycontact 17 28 17 28 1 b
rlabel pdiffusion 14 37 14 37 1 d1s2
rlabel metal1 41 25 41 25 3 out
rlabel metal1 24 22 24 22 5 toInv
rlabel polycontact 34 22 34 22 1 inv
<< end >>
