magic
tech scmos
timestamp 1635707612
<< nwell >>
rect -11 2 24 13
<< polysilicon >>
rect -5 10 -3 12
rect 5 10 7 12
rect 15 10 17 12
rect -5 -2 -3 4
rect -4 -6 -3 -2
rect 5 -5 7 4
rect 15 -5 17 4
rect -5 -10 -3 -6
rect 6 -9 7 -5
rect 16 -9 17 -5
rect 5 -10 7 -9
rect 15 -10 17 -9
rect -5 -21 -3 -19
rect 5 -21 7 -19
rect 15 -21 17 -19
<< ndiffusion >>
rect -10 -13 -5 -10
rect -7 -17 -5 -13
rect -10 -19 -5 -17
rect -3 -19 5 -10
rect 7 -19 15 -10
rect 17 -13 23 -10
rect 17 -17 19 -13
rect 17 -19 23 -17
<< pdiffusion >>
rect -10 9 -5 10
rect -7 5 -5 9
rect -10 4 -5 5
rect -3 9 5 10
rect -3 5 -1 9
rect 3 5 5 9
rect -3 4 5 5
rect 7 9 15 10
rect 7 5 9 9
rect 13 5 15 9
rect 7 4 15 5
rect 17 9 23 10
rect 17 5 19 9
rect 17 4 23 5
<< metal1 >>
rect -11 16 1 18
rect 5 16 12 18
rect -11 15 12 16
rect -11 9 -8 15
rect 9 9 12 15
rect 0 1 3 5
rect 20 1 23 5
rect 0 -2 23 1
rect 20 -13 23 -2
rect -11 -23 -8 -17
rect -11 -24 9 -23
rect -11 -26 4 -24
rect 8 -26 9 -24
<< ntransistor >>
rect -5 -19 -3 -10
rect 5 -19 7 -10
rect 15 -19 17 -10
<< ptransistor >>
rect -5 4 -3 10
rect 5 4 7 10
rect 15 4 17 10
<< polycontact >>
rect -8 -6 -4 -2
rect 2 -9 6 -5
rect 12 -9 16 -5
<< ndcontact >>
rect -11 -17 -7 -13
rect 19 -17 23 -13
<< pdcontact >>
rect -11 5 -7 9
rect -1 5 3 9
rect 9 5 13 9
rect 19 5 23 9
<< psubstratepcontact >>
rect 4 -28 8 -24
<< nsubstratencontact >>
rect 1 16 5 20
<< labels >>
rlabel metal1 -3 -25 -3 -25 1 vss
rlabel metal1 -6 16 -6 16 1 vdd
rlabel metal1 21 -1 21 -1 1 out
rlabel polycontact -6 -4 -6 -4 1 C
rlabel polycontact 4 -7 4 -7 1 B
rlabel polycontact 14 -7 14 -7 1 A
rlabel ndiffusion 1 -15 1 -15 1 s2d3
rlabel ndiffusion 11 -15 11 -15 1 s1d2
<< end >>
