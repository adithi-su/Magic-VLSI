magic
tech scmos
timestamp 1636302090
<< nwell >>
rect 68 86 100 103
rect 6 63 38 80
rect 126 76 158 93
rect 248 86 280 103
rect 186 63 218 80
rect 306 76 338 93
rect 68 37 100 54
rect 136 32 156 48
rect 248 37 280 54
rect 316 32 336 48
rect 348 40 397 55
<< polysilicon >>
rect 73 94 75 96
rect 93 94 95 96
rect 253 94 255 96
rect 273 94 275 96
rect 73 86 75 88
rect 74 82 75 86
rect 11 71 13 73
rect 31 71 33 73
rect 73 71 75 82
rect 93 79 95 88
rect 253 86 255 88
rect 131 84 133 86
rect 151 84 153 86
rect 94 75 95 79
rect 254 82 255 86
rect 131 76 133 78
rect 93 71 95 75
rect 132 72 133 76
rect 73 66 75 68
rect 93 66 95 68
rect 11 63 13 65
rect 12 59 13 63
rect 11 48 13 59
rect 31 56 33 65
rect 131 61 133 72
rect 151 69 153 78
rect 191 71 193 73
rect 211 71 213 73
rect 152 65 153 69
rect 253 71 255 82
rect 273 79 275 88
rect 311 84 313 86
rect 331 84 333 86
rect 274 75 275 79
rect 311 76 313 78
rect 273 71 275 75
rect 312 72 313 76
rect 253 66 255 68
rect 273 66 275 68
rect 151 61 153 65
rect 191 63 193 65
rect 192 59 193 63
rect 131 56 133 58
rect 151 56 153 58
rect 32 52 33 56
rect 31 48 33 52
rect 73 45 75 47
rect 93 45 95 47
rect 11 43 13 45
rect 31 43 33 45
rect 191 48 193 59
rect 211 56 213 65
rect 311 61 313 72
rect 331 69 333 78
rect 332 65 333 69
rect 331 61 333 65
rect 311 56 313 58
rect 331 56 333 58
rect 212 52 213 56
rect 211 48 213 52
rect 253 45 255 47
rect 273 45 275 47
rect 191 43 193 45
rect 211 43 213 45
rect 144 39 146 41
rect 353 47 355 49
rect 369 47 371 49
rect 389 47 391 49
rect 324 39 326 41
rect 73 37 75 39
rect 74 33 75 37
rect 73 22 75 33
rect 93 30 95 39
rect 253 37 255 39
rect 254 33 255 37
rect 144 30 146 33
rect 94 26 95 30
rect 93 22 95 26
rect 144 22 146 26
rect 73 17 75 19
rect 93 17 95 19
rect 144 17 146 19
rect 253 22 255 33
rect 273 30 275 39
rect 324 30 326 33
rect 274 26 275 30
rect 353 29 355 41
rect 369 38 371 41
rect 370 34 371 38
rect 273 22 275 26
rect 324 22 326 26
rect 354 25 355 29
rect 253 17 255 19
rect 273 17 275 19
rect 324 17 326 19
rect 353 21 355 25
rect 369 21 371 34
rect 389 29 391 41
rect 389 22 391 25
rect 353 16 355 18
rect 369 16 371 18
rect 389 16 391 18
<< ndiffusion >>
rect 72 68 73 71
rect 75 68 93 71
rect 95 68 96 71
rect 252 68 253 71
rect 255 68 273 71
rect 275 68 276 71
rect 130 58 131 61
rect 133 58 151 61
rect 153 58 154 61
rect 10 45 11 48
rect 13 45 31 48
rect 33 45 34 48
rect 310 58 311 61
rect 313 58 331 61
rect 333 58 334 61
rect 190 45 191 48
rect 193 45 211 48
rect 213 45 214 48
rect 72 19 73 22
rect 75 19 93 22
rect 95 19 96 22
rect 142 19 144 22
rect 146 19 148 22
rect 252 19 253 22
rect 255 19 273 22
rect 275 19 276 22
rect 322 19 324 22
rect 326 19 328 22
rect 352 18 353 21
rect 355 18 356 21
rect 368 18 369 21
rect 371 18 372 21
rect 387 18 389 22
rect 391 18 393 22
<< pdiffusion >>
rect 70 93 73 94
rect 72 89 73 93
rect 70 88 73 89
rect 75 93 78 94
rect 90 93 93 94
rect 75 89 76 93
rect 92 89 93 93
rect 75 88 78 89
rect 90 88 93 89
rect 95 93 98 94
rect 250 93 253 94
rect 95 89 96 93
rect 252 89 253 93
rect 95 88 98 89
rect 250 88 253 89
rect 255 93 258 94
rect 270 93 273 94
rect 255 89 256 93
rect 272 89 273 93
rect 255 88 258 89
rect 270 88 273 89
rect 275 93 278 94
rect 275 89 276 93
rect 275 88 278 89
rect 8 70 11 71
rect 10 66 11 70
rect 8 65 11 66
rect 13 70 16 71
rect 28 70 31 71
rect 13 66 14 70
rect 30 66 31 70
rect 13 65 16 66
rect 28 65 31 66
rect 33 70 36 71
rect 33 66 34 70
rect 128 83 131 84
rect 130 79 131 83
rect 128 78 131 79
rect 133 83 136 84
rect 148 83 151 84
rect 133 79 134 83
rect 150 79 151 83
rect 133 78 136 79
rect 148 78 151 79
rect 153 83 156 84
rect 153 79 154 83
rect 153 78 156 79
rect 33 65 36 66
rect 188 70 191 71
rect 190 66 191 70
rect 188 65 191 66
rect 193 70 196 71
rect 208 70 211 71
rect 193 66 194 70
rect 210 66 211 70
rect 193 65 196 66
rect 208 65 211 66
rect 213 70 216 71
rect 213 66 214 70
rect 308 83 311 84
rect 310 79 311 83
rect 308 78 311 79
rect 313 83 316 84
rect 328 83 331 84
rect 313 79 314 83
rect 330 79 331 83
rect 313 78 316 79
rect 328 78 331 79
rect 333 83 336 84
rect 333 79 334 83
rect 333 78 336 79
rect 213 65 216 66
rect 70 44 73 45
rect 72 40 73 44
rect 70 39 73 40
rect 75 44 78 45
rect 90 44 93 45
rect 75 40 76 44
rect 92 40 93 44
rect 75 39 78 40
rect 90 39 93 40
rect 95 44 98 45
rect 95 40 96 44
rect 250 44 253 45
rect 95 39 98 40
rect 252 40 253 44
rect 250 39 253 40
rect 255 44 258 45
rect 270 44 273 45
rect 255 40 256 44
rect 272 40 273 44
rect 255 39 258 40
rect 270 39 273 40
rect 275 44 278 45
rect 350 46 353 47
rect 275 40 276 44
rect 352 42 353 46
rect 350 41 353 42
rect 355 41 369 47
rect 371 46 375 47
rect 384 46 389 47
rect 371 42 372 46
rect 387 42 389 46
rect 371 41 375 42
rect 384 41 389 42
rect 391 46 396 47
rect 391 42 393 46
rect 391 41 396 42
rect 275 39 278 40
rect 141 38 144 39
rect 143 34 144 38
rect 141 33 144 34
rect 146 38 150 39
rect 146 34 147 38
rect 146 33 150 34
rect 321 38 324 39
rect 323 34 324 38
rect 321 33 324 34
rect 326 38 330 39
rect 326 34 327 38
rect 326 33 330 34
<< metal1 >>
rect 20 99 60 102
rect 64 99 68 102
rect 72 99 88 102
rect 92 99 126 102
rect 130 99 196 102
rect 200 99 240 102
rect 244 99 248 102
rect 252 99 268 102
rect 272 99 306 102
rect 310 99 345 102
rect 69 93 72 99
rect 88 93 91 99
rect 127 93 130 99
rect 130 89 146 92
rect 77 86 80 89
rect 97 86 100 89
rect 0 83 70 86
rect 0 63 3 83
rect 77 83 100 86
rect 127 83 130 89
rect 146 83 149 89
rect 10 76 16 79
rect 20 76 26 79
rect 7 70 10 76
rect 26 70 29 76
rect 44 75 90 78
rect 97 76 100 83
rect 135 76 138 79
rect 155 76 158 79
rect 15 63 18 66
rect 35 63 38 66
rect 44 63 47 75
rect 97 73 128 76
rect 97 72 100 73
rect 135 73 158 76
rect 155 72 158 73
rect 68 64 71 68
rect 103 65 148 68
rect 155 68 156 72
rect 0 60 8 63
rect 15 60 47 63
rect 57 60 68 63
rect 0 53 28 56
rect 0 30 3 53
rect 35 49 38 60
rect 6 37 9 45
rect 44 38 47 60
rect 64 50 68 53
rect 72 50 88 53
rect 69 44 72 50
rect 88 44 91 50
rect 77 37 80 40
rect 97 37 100 40
rect 103 37 106 65
rect 155 62 158 68
rect 48 34 70 37
rect 77 34 106 37
rect 0 27 90 30
rect 97 23 100 34
rect 68 15 71 19
rect 126 15 129 58
rect 139 44 150 45
rect 164 47 167 99
rect 249 93 252 99
rect 268 93 271 99
rect 307 93 310 99
rect 310 89 326 92
rect 257 86 260 89
rect 277 86 280 89
rect 180 83 250 86
rect 180 63 183 83
rect 257 83 280 86
rect 307 83 310 89
rect 326 83 329 89
rect 190 76 196 79
rect 200 76 206 79
rect 187 70 190 76
rect 206 70 209 76
rect 224 75 270 78
rect 277 76 280 83
rect 315 76 318 79
rect 335 76 338 79
rect 195 63 198 66
rect 215 63 218 66
rect 224 63 227 75
rect 277 73 308 76
rect 277 72 280 73
rect 315 73 338 76
rect 248 64 251 68
rect 283 65 328 68
rect 180 60 188 63
rect 195 60 227 63
rect 237 60 248 63
rect 154 44 167 47
rect 180 53 208 56
rect 180 45 183 53
rect 215 49 218 60
rect 139 42 153 44
rect 139 38 142 42
rect 182 40 183 45
rect 151 34 153 38
rect 136 26 142 29
rect 150 29 153 34
rect 180 30 183 40
rect 186 37 189 45
rect 224 38 227 60
rect 244 50 248 53
rect 252 50 268 53
rect 249 44 252 50
rect 268 44 271 50
rect 257 37 260 40
rect 277 37 280 40
rect 283 37 286 65
rect 335 62 338 73
rect 228 34 250 37
rect 257 34 286 37
rect 150 25 151 29
rect 180 27 270 30
rect 150 22 153 25
rect 277 23 280 34
rect 152 18 153 22
rect 138 15 141 18
rect 248 15 251 19
rect 306 15 309 58
rect 342 55 345 99
rect 342 52 348 55
rect 319 44 330 45
rect 342 47 345 52
rect 334 44 345 47
rect 352 52 383 55
rect 348 46 351 51
rect 383 46 386 51
rect 319 42 333 44
rect 319 38 322 42
rect 331 37 333 38
rect 331 34 366 37
rect 316 26 322 29
rect 330 22 333 34
rect 343 25 350 28
rect 373 28 376 42
rect 357 25 387 28
rect 357 22 360 25
rect 373 22 376 25
rect 394 22 397 42
rect 332 18 333 22
rect 318 15 321 18
rect 348 15 351 18
rect 364 15 367 18
rect 384 15 387 18
rect 10 12 28 15
rect 32 12 54 15
rect 58 12 68 15
rect 72 12 96 15
rect 100 12 125 15
rect 129 14 186 15
rect 129 12 148 14
rect 152 12 186 14
rect 190 12 208 15
rect 212 12 234 15
rect 238 12 248 15
rect 252 12 276 15
rect 280 12 305 15
rect 309 14 387 15
rect 309 12 328 14
rect 332 12 360 14
rect 364 12 387 14
rect 166 0 339 3
<< metal2 >>
rect 17 80 20 99
rect 6 15 9 33
rect 45 7 48 34
rect 53 15 56 60
rect 61 54 64 99
rect 197 80 200 99
rect 160 68 175 71
rect 172 45 175 68
rect 172 42 177 45
rect 182 42 183 45
rect 53 12 54 15
rect 132 7 135 26
rect 155 26 165 29
rect 45 4 135 7
rect 162 4 165 26
rect 186 15 189 33
rect 225 7 228 34
rect 233 15 236 60
rect 241 54 244 99
rect 233 12 234 15
rect 312 7 315 26
rect 225 4 315 7
rect 340 4 343 25
<< ntransistor >>
rect 73 68 75 71
rect 93 68 95 71
rect 253 68 255 71
rect 273 68 275 71
rect 131 58 133 61
rect 151 58 153 61
rect 11 45 13 48
rect 31 45 33 48
rect 311 58 313 61
rect 331 58 333 61
rect 191 45 193 48
rect 211 45 213 48
rect 73 19 75 22
rect 93 19 95 22
rect 144 19 146 22
rect 253 19 255 22
rect 273 19 275 22
rect 324 19 326 22
rect 353 18 355 21
rect 369 18 371 21
rect 389 18 391 22
<< ptransistor >>
rect 73 88 75 94
rect 93 88 95 94
rect 253 88 255 94
rect 273 88 275 94
rect 11 65 13 71
rect 31 65 33 71
rect 131 78 133 84
rect 151 78 153 84
rect 191 65 193 71
rect 211 65 213 71
rect 311 78 313 84
rect 331 78 333 84
rect 73 39 75 45
rect 93 39 95 45
rect 253 39 255 45
rect 273 39 275 45
rect 353 41 355 47
rect 369 41 371 47
rect 389 41 391 47
rect 144 33 146 39
rect 324 33 326 39
<< polycontact >>
rect 70 82 74 86
rect 90 75 94 79
rect 250 82 254 86
rect 128 72 132 76
rect 8 59 12 63
rect 148 65 152 69
rect 270 75 274 79
rect 308 72 312 76
rect 188 59 192 63
rect 28 52 32 56
rect 328 65 332 69
rect 208 52 212 56
rect 70 33 74 37
rect 250 33 254 37
rect 90 26 94 30
rect 142 26 146 30
rect 270 26 274 30
rect 322 26 326 30
rect 366 34 370 38
rect 350 25 354 29
rect 387 25 391 29
<< ndcontact >>
rect 68 68 72 72
rect 96 68 100 72
rect 6 45 10 49
rect 126 58 130 62
rect 248 68 252 72
rect 276 68 280 72
rect 154 58 158 62
rect 34 45 38 49
rect 186 45 190 49
rect 306 58 310 62
rect 334 58 338 62
rect 214 45 218 49
rect 68 19 72 23
rect 96 19 100 23
rect 138 18 142 22
rect 148 18 152 22
rect 248 19 252 23
rect 276 19 280 23
rect 318 18 322 22
rect 328 18 332 22
rect 348 18 352 22
rect 356 18 360 22
rect 364 18 368 22
rect 372 18 376 22
rect 383 18 387 22
rect 393 18 397 22
<< pdcontact >>
rect 68 89 72 93
rect 76 89 80 93
rect 88 89 92 93
rect 96 89 100 93
rect 248 89 252 93
rect 256 89 260 93
rect 268 89 272 93
rect 276 89 280 93
rect 6 66 10 70
rect 14 66 18 70
rect 26 66 30 70
rect 34 66 38 70
rect 126 79 130 83
rect 134 79 138 83
rect 146 79 150 83
rect 154 79 158 83
rect 186 66 190 70
rect 194 66 198 70
rect 206 66 210 70
rect 214 66 218 70
rect 306 79 310 83
rect 314 79 318 83
rect 326 79 330 83
rect 334 79 338 83
rect 68 40 72 44
rect 76 40 80 44
rect 88 40 92 44
rect 96 40 100 44
rect 248 40 252 44
rect 256 40 260 44
rect 268 40 272 44
rect 276 40 280 44
rect 348 42 352 46
rect 372 42 376 46
rect 383 42 387 46
rect 393 42 397 46
rect 139 34 143 38
rect 147 34 151 38
rect 319 34 323 38
rect 327 34 331 38
<< m2contact >>
rect 16 99 20 103
rect 60 99 64 103
rect 196 99 200 103
rect 240 99 244 103
rect 16 76 20 80
rect 156 68 160 72
rect 53 60 57 64
rect 60 50 64 54
rect 6 33 10 37
rect 44 34 48 38
rect 196 76 200 80
rect 233 60 237 64
rect 177 40 182 45
rect 132 26 136 30
rect 240 50 244 54
rect 186 33 190 37
rect 224 34 228 38
rect 151 25 155 29
rect 312 26 316 30
rect 339 25 343 29
rect 6 11 10 15
rect 54 11 58 15
rect 186 11 190 15
rect 234 11 238 15
rect 162 0 166 4
rect 339 0 343 4
<< psubstratepcontact >>
rect 68 60 72 64
rect 248 60 252 64
rect 28 11 32 15
rect 68 11 72 15
rect 96 11 100 15
rect 125 11 129 15
rect 148 10 152 14
rect 208 11 212 15
rect 248 11 252 15
rect 276 11 280 15
rect 305 11 309 15
rect 328 10 332 14
rect 360 10 364 14
<< nsubstratencontact >>
rect 68 99 72 103
rect 88 99 92 103
rect 126 99 130 103
rect 248 99 252 103
rect 268 99 272 103
rect 306 99 310 103
rect 126 89 130 93
rect 146 89 150 93
rect 306 89 310 93
rect 326 89 330 93
rect 6 76 10 80
rect 26 76 30 80
rect 186 76 190 80
rect 206 76 210 80
rect 68 50 72 54
rect 88 50 92 54
rect 150 44 154 48
rect 248 50 252 54
rect 268 50 272 54
rect 348 51 352 55
rect 383 51 387 55
rect 330 44 334 48
<< labels >>
rlabel polycontact 252 84 252 84 1 A
rlabel polycontact 190 61 190 61 1 A
rlabel polycontact 272 28 272 28 1 B
rlabel polycontact 210 54 210 54 1 B
rlabel metal1 181 28 181 28 1 B
rlabel metal1 218 13 218 13 1 Gnd
rlabel metal1 221 100 221 100 1 Vdd
rlabel metal1 336 74 336 74 1 sum
rlabel metal1 38 13 38 13 1 Gnd
rlabel metal1 41 100 41 100 1 Vdd
rlabel metal1 156 74 156 74 1 sum1
rlabel polycontact 92 28 92 28 1 B1
rlabel polycontact 72 84 72 84 1 A1
rlabel polycontact 30 54 30 54 1 B1
rlabel polycontact 10 61 10 61 1 A1
rlabel metal1 1 28 1 28 1 B1
rlabel metal1 1 84 1 84 1 A1
rlabel metal1 181 84 181 84 3 C_in
rlabel metal1 330 1 330 1 1 carry2
rlabel metal1 355 13 355 13 3 Gnd
rlabel metal1 396 31 396 31 1 C_out
rlabel metal1 366 53 366 53 1 Vdd
rlabel metal1 331 27 331 27 1 carry1
<< end >>
