magic
tech scmos
timestamp 1635704755
<< nwell >>
rect -14 7 12 20
<< polysilicon >>
rect -7 16 -5 18
rect 4 16 6 18
rect -7 4 -5 10
rect 4 6 6 10
rect -6 0 -5 4
rect 5 2 6 6
rect -7 -8 -5 0
rect 4 -8 6 2
rect -7 -17 -5 -14
rect 4 -17 6 -14
<< ndiffusion >>
rect -12 -9 -7 -8
rect -9 -13 -7 -9
rect -12 -14 -7 -13
rect -5 -9 4 -8
rect -5 -13 -2 -9
rect 2 -13 4 -9
rect -5 -14 4 -13
rect 6 -9 10 -8
rect 6 -13 8 -9
rect 6 -14 10 -13
<< pdiffusion >>
rect -12 15 -7 16
rect -9 11 -7 15
rect -12 10 -7 11
rect -5 10 4 16
rect 6 15 10 16
rect 6 11 8 15
rect 6 10 10 11
<< metal1 >>
rect -13 22 0 25
rect 4 22 8 25
rect -13 15 -10 22
rect 9 -1 12 11
rect -2 -4 12 -1
rect -2 -9 1 -4
rect -12 -19 -9 -13
rect 9 -19 12 -13
rect -12 -20 12 -19
rect -12 -22 -1 -20
rect 3 -22 12 -20
<< ntransistor >>
rect -7 -14 -5 -8
rect 4 -14 6 -8
<< ptransistor >>
rect -7 10 -5 16
rect 4 10 6 16
<< polycontact >>
rect -10 0 -6 4
rect 1 2 5 6
<< ndcontact >>
rect -13 -13 -9 -9
rect -2 -13 2 -9
rect 8 -13 12 -9
<< pdcontact >>
rect -13 11 -9 15
rect 8 11 12 15
<< psubstratepcontact >>
rect -1 -24 3 -20
<< nsubstratencontact >>
rect 0 22 4 26
<< labels >>
rlabel metal1 -5 23 -5 23 1 vdd
rlabel metal1 -6 -21 -6 -21 1 vss
rlabel polycontact -8 2 -8 2 1 a
rlabel polycontact 3 4 3 4 1 b
rlabel metal1 11 0 11 0 7 out
rlabel pdiffusion 0 13 0 13 1 d1s2
<< end >>
