magic
tech scmos
timestamp 1635798489
<< nwell >>
rect 31 49 57 60
rect 0 22 20 38
rect 27 -5 53 6
<< polysilicon >>
rect 36 57 38 60
rect 49 57 51 60
rect 36 42 38 51
rect 37 38 38 42
rect 49 39 51 51
rect 36 31 38 38
rect 50 35 51 39
rect 49 31 51 35
rect 8 29 10 31
rect 36 23 38 25
rect 49 23 51 25
rect 8 19 10 23
rect 9 15 10 19
rect 8 12 10 15
rect 8 7 10 9
rect 32 3 34 6
rect 45 3 47 6
rect 32 -12 34 -3
rect 33 -16 34 -12
rect 45 -15 47 -3
rect 32 -23 34 -16
rect 46 -19 47 -15
rect 45 -23 47 -19
rect 32 -31 34 -29
rect 45 -31 47 -29
<< ndiffusion >>
rect 32 30 36 31
rect 34 26 36 30
rect 32 25 36 26
rect 38 25 49 31
rect 51 30 55 31
rect 51 26 53 30
rect 51 25 55 26
rect 6 9 8 12
rect 10 9 12 12
rect 28 -24 32 -23
rect 30 -28 32 -24
rect 28 -29 32 -28
rect 34 -29 45 -23
rect 47 -24 51 -23
rect 47 -28 49 -24
rect 47 -29 51 -28
<< pdiffusion >>
rect 32 56 36 57
rect 34 52 36 56
rect 32 51 36 52
rect 38 56 49 57
rect 38 52 41 56
rect 45 52 49 56
rect 38 51 49 52
rect 51 56 55 57
rect 51 52 53 56
rect 51 51 55 52
rect 5 28 8 29
rect 7 24 8 28
rect 5 23 8 24
rect 10 28 14 29
rect 10 24 11 28
rect 10 23 14 24
rect 28 2 32 3
rect 30 -2 32 2
rect 28 -3 32 -2
rect 34 2 45 3
rect 34 -2 37 2
rect 41 -2 45 2
rect 34 -3 45 -2
rect 47 2 51 3
rect 47 -2 49 2
rect 47 -3 51 -2
<< metal1 >>
rect 33 63 45 65
rect 49 63 57 65
rect 33 62 57 63
rect 30 56 33 62
rect 54 56 57 62
rect 42 47 45 52
rect 42 44 54 47
rect 22 38 33 41
rect 3 33 6 35
rect 10 33 14 35
rect 3 32 17 33
rect 3 28 6 32
rect 15 24 17 28
rect 14 20 17 24
rect 22 20 25 38
rect 54 30 57 43
rect -4 15 5 18
rect 14 17 25 20
rect 30 22 33 26
rect 30 20 60 22
rect -4 -13 -1 15
rect 14 12 17 17
rect 34 19 60 20
rect 16 8 17 12
rect 2 5 5 8
rect 29 9 41 11
rect 45 9 53 11
rect 29 8 53 9
rect 2 4 15 5
rect 2 2 5 4
rect 9 2 12 4
rect 26 2 29 7
rect 50 2 53 8
rect 38 -7 41 -2
rect 38 -10 50 -7
rect -4 -16 29 -13
rect 50 -24 53 -11
rect 26 -32 29 -28
rect 57 -32 60 19
rect 10 -33 60 -32
rect 10 -35 38 -33
rect 42 -35 60 -33
<< metal2 >>
rect 7 62 29 65
rect 7 37 10 62
rect 26 11 29 62
rect 58 44 73 47
rect 48 35 65 38
rect 6 -32 9 0
rect 62 -7 65 35
rect 54 -10 65 -7
rect 70 -16 73 44
rect 44 -19 73 -16
<< ntransistor >>
rect 36 25 38 31
rect 49 25 51 31
rect 8 9 10 12
rect 32 -29 34 -23
rect 45 -29 47 -23
<< ptransistor >>
rect 36 51 38 57
rect 49 51 51 57
rect 8 23 10 29
rect 32 -3 34 3
rect 45 -3 47 3
<< polycontact >>
rect 33 38 37 42
rect 46 35 50 39
rect 5 15 9 19
rect 29 -16 33 -12
rect 42 -19 46 -15
<< ndcontact >>
rect 30 26 34 30
rect 53 26 57 30
rect 2 8 6 12
rect 12 8 16 12
rect 26 -28 30 -24
rect 49 -28 53 -24
<< pdcontact >>
rect 30 52 34 56
rect 41 52 45 56
rect 53 52 57 56
rect 3 24 7 28
rect 11 24 15 28
rect 26 -2 30 2
rect 37 -2 41 2
rect 49 -2 53 2
<< m2contact >>
rect 29 62 33 66
rect 54 43 58 47
rect 6 33 10 37
rect 25 7 29 11
rect 5 0 9 4
rect 50 -11 54 -7
rect 6 -36 10 -32
<< psubstratepcontact >>
rect 30 16 34 20
rect 12 0 16 4
rect 38 -37 42 -33
<< nsubstratencontact >>
rect 45 63 49 67
rect 14 33 18 37
rect 41 9 45 13
<< labels >>
rlabel metal1 15 15 15 15 1 D_bar
rlabel polycontact 31 -14 31 -14 1 D
rlabel metal1 28 -34 28 -34 1 vss
rlabel metal1 51 -13 51 -13 3 Q_bar
rlabel metal1 55 40 55 40 3 Q
rlabel polycontact 35 40 35 40 1 D_bar
rlabel metal1 36 64 36 64 5 vdd
rlabel polycontact 7 17 7 17 1 in
<< end >>
