magic
tech scmos
timestamp 1635706314
<< nwell >>
rect -12 5 14 16
<< polysilicon >>
rect -7 13 -5 16
rect 6 13 8 16
rect -7 -2 -5 7
rect -6 -6 -5 -2
rect 6 -5 8 7
rect -7 -13 -5 -6
rect 7 -9 8 -5
rect 6 -13 8 -9
rect -7 -21 -5 -19
rect 6 -21 8 -19
<< ndiffusion >>
rect -11 -14 -7 -13
rect -9 -18 -7 -14
rect -11 -19 -7 -18
rect -5 -19 6 -13
rect 8 -14 12 -13
rect 8 -18 10 -14
rect 8 -19 12 -18
<< pdiffusion >>
rect -11 12 -7 13
rect -9 8 -7 12
rect -11 7 -7 8
rect -5 12 6 13
rect -5 8 -2 12
rect 2 8 6 12
rect -5 7 6 8
rect 8 12 12 13
rect 8 8 10 12
rect 8 7 12 8
<< metal1 >>
rect -13 19 2 21
rect 6 19 14 21
rect -13 18 14 19
rect -13 12 -10 18
rect 11 12 14 18
rect -1 3 2 8
rect -1 0 14 3
rect 11 -14 14 0
rect -13 -22 -10 -18
rect -13 -23 3 -22
rect -13 -25 -1 -23
<< ntransistor >>
rect -7 -19 -5 -13
rect 6 -19 8 -13
<< ptransistor >>
rect -7 7 -5 13
rect 6 7 8 13
<< polycontact >>
rect -10 -6 -6 -2
rect 3 -9 7 -5
<< ndcontact >>
rect -13 -18 -9 -14
rect 10 -18 14 -14
<< pdcontact >>
rect -13 8 -9 12
rect -2 8 2 12
rect 10 8 14 12
<< psubstratepcontact >>
rect -1 -27 3 -23
<< nsubstratencontact >>
rect 2 19 6 23
<< labels >>
rlabel polycontact -8 -4 -8 -4 1 b
rlabel polycontact 5 -7 5 -7 1 a
rlabel metal1 -11 -24 -11 -24 1 vss
rlabel metal1 12 -3 12 -3 3 out
rlabel metal1 -7 20 -7 20 5 vdd
rlabel ndiffusion 1 -16 1 -16 1 s1d2
<< end >>
