* SPICE3 file created from and2.ext - technology: scmos

.option scale=1u

M1000 vdd a inv vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 inv a s1d2 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 inv b vdd vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out inv vdd vdd pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 out inv inv Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 s1d2 b inv Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out Gnd 2.58fF
C1 inv Gnd 16.34fF
C2 a Gnd 6.19fF
C3 b Gnd 6.19fF
