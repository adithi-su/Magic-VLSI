magic
tech scmos
timestamp 1635711265
<< nwell >>
rect -1 32 48 49
<< polysilicon >>
rect 6 40 8 43
rect 19 40 21 43
rect 37 40 39 43
rect 6 25 8 34
rect 7 21 8 25
rect 19 22 21 34
rect 37 30 39 34
rect 38 26 39 30
rect 6 14 8 21
rect 20 18 21 22
rect 19 14 21 18
rect 37 14 39 26
rect 6 6 8 8
rect 19 6 21 8
rect 37 6 39 8
<< ndiffusion >>
rect 2 13 6 14
rect 4 9 6 13
rect 2 8 6 9
rect 8 8 19 14
rect 21 13 37 14
rect 21 9 23 13
rect 27 9 30 13
rect 34 9 37 13
rect 21 8 37 9
rect 39 13 44 14
rect 39 9 41 13
rect 39 8 44 9
<< pdiffusion >>
rect 2 39 6 40
rect 4 35 6 39
rect 2 34 6 35
rect 8 39 19 40
rect 8 35 11 39
rect 15 35 19 39
rect 8 34 19 35
rect 21 39 37 40
rect 21 35 28 39
rect 32 35 37 39
rect 21 34 37 35
rect 39 39 43 40
rect 39 35 41 39
rect 39 34 43 35
<< metal1 >>
rect 0 46 15 48
rect 19 46 31 48
rect 0 45 31 46
rect 0 39 3 45
rect 28 39 31 45
rect 12 30 15 35
rect 12 27 34 30
rect 24 13 27 27
rect 42 13 45 35
rect 0 5 3 9
rect 30 5 33 9
rect 0 4 33 5
rect 0 2 12 4
rect 16 2 33 4
<< ntransistor >>
rect 6 8 8 14
rect 19 8 21 14
rect 37 8 39 14
<< ptransistor >>
rect 6 34 8 40
rect 19 34 21 40
rect 37 34 39 40
<< polycontact >>
rect 3 21 7 25
rect 34 26 38 30
rect 16 18 20 22
<< ndcontact >>
rect 0 9 4 13
rect 23 9 27 13
rect 30 9 34 13
rect 41 9 45 13
<< pdcontact >>
rect 0 35 4 39
rect 11 35 15 39
rect 28 35 32 39
rect 41 35 45 39
<< psubstratepcontact >>
rect 12 0 16 4
<< nsubstratencontact >>
rect 15 46 19 50
<< labels >>
rlabel polycontact 5 23 5 23 1 b
rlabel polycontact 18 20 18 20 1 a
rlabel metal1 2 3 2 3 1 vss
rlabel metal1 6 47 6 47 5 vdd
rlabel ndiffusion 14 11 14 11 1 s1d2
rlabel metal1 44 24 44 24 7 out
rlabel metal1 26 28 26 28 1 toInv
rlabel polycontact 36 28 36 28 1 inv
<< end >>
