magic
tech scmos
timestamp 1635719768
<< nwell >>
rect -16 1 37 16
<< polysilicon >>
rect -11 10 -9 12
rect 0 10 2 12
rect 17 10 19 12
rect 27 10 29 12
rect -11 -6 -9 2
rect 0 -6 2 2
rect 17 -2 19 2
rect 18 -6 19 -2
rect -10 -10 -9 -6
rect 1 -10 2 -6
rect -11 -20 -9 -10
rect 0 -20 2 -10
rect 17 -20 19 -6
rect 27 -13 29 2
rect 27 -17 28 -13
rect 27 -20 29 -17
rect -11 -27 -9 -25
rect 0 -27 2 -25
rect 17 -27 19 -25
rect 27 -27 29 -25
<< ndiffusion >>
rect -15 -21 -11 -20
rect -13 -25 -11 -21
rect -9 -25 0 -20
rect 2 -21 17 -20
rect 2 -25 7 -21
rect 11 -25 17 -21
rect 19 -25 27 -20
rect 29 -21 35 -20
rect 29 -25 31 -21
<< pdiffusion >>
rect -14 7 -11 10
rect -12 3 -11 7
rect -14 2 -11 3
rect -9 7 0 10
rect -9 3 -6 7
rect -2 3 0 7
rect -9 2 0 3
rect 2 7 17 10
rect 2 3 4 7
rect 8 3 11 7
rect 15 3 17 7
rect 2 2 17 3
rect 19 7 27 10
rect 19 3 21 7
rect 25 3 27 7
rect 19 2 27 3
rect 29 7 36 10
rect 29 3 31 7
rect 35 3 36 7
rect 29 2 36 3
<< metal1 >>
rect -12 14 7 16
rect -16 13 7 14
rect -16 7 -13 13
rect 4 7 7 13
rect 22 -9 25 3
rect 8 -12 25 -9
rect 8 -21 11 -12
rect -16 -29 -13 -25
rect 31 -29 34 -25
rect -16 -32 7 -29
rect 11 -32 34 -29
<< metal2 >>
rect -5 19 34 22
rect -5 4 -2 19
rect 11 4 14 19
rect 31 4 34 19
<< ntransistor >>
rect -11 -25 -9 -20
rect 0 -25 2 -20
rect 17 -25 19 -20
rect 27 -25 29 -20
<< ptransistor >>
rect -11 2 -9 10
rect 0 2 2 10
rect 17 2 19 10
rect 27 2 29 10
<< polycontact >>
rect 14 -6 18 -2
rect -14 -10 -10 -6
rect -3 -10 1 -6
rect 28 -17 32 -13
<< ndcontact >>
rect -17 -25 -13 -21
rect 7 -25 11 -21
rect 31 -25 35 -21
<< pdcontact >>
rect -16 3 -12 7
rect -6 3 -2 7
rect 4 3 8 7
rect 11 3 15 7
rect 21 3 25 7
rect 31 3 35 7
<< psubstratepcontact >>
rect 7 -33 11 -29
<< nsubstratencontact >>
rect -16 14 -12 18
<< labels >>
rlabel metal1 23 -10 23 -10 3 out
rlabel metal1 -7 -31 -7 -31 1 vss
rlabel polycontact -12 -8 -12 -8 1 B
rlabel polycontact -1 -8 -1 -8 1 A
rlabel polycontact 16 -4 16 -4 1 C
rlabel polycontact 30 -15 30 -15 1 D
rlabel metal1 -10 14 -10 14 1 vdd
<< end >>
