* SPICE3 file created from nand2.ext - technology: scmos

.option scale=1u

M1000 out b vdd w_n12_5# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 s1d2 b vss Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 vdd a out w_n12_5# pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out a s1d2 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vss Gnd 2.40fF
C1 out Gnd 4.04fF
C2 a Gnd 6.35fF
C3 b Gnd 6.35fF
C4 vdd Gnd 4.18fF
